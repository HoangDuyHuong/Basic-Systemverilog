package math_pkg;

function int plus (int a, int b);
	plus = a+b;
endfunction

function int minus (int a, int b);
	minus = a-b;
endfunction

endpackage

